//Alot of things